


 






// file: ibert_7series_gtp_3750.v
//////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2012.3
//  \   \         Application : IBERT 7Series 
//  /   /         Filename : example_ibert_7series_gtp_3750
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\
//
//
// Module example_ibert_7series_gtp_3750
// Generated by Xilinx IBERT_7S 
//////////////////////////////////////////////////////////////////////////////


`define C_NUM_QUADS 1
`define C_REFCLKS_USED 1
module example_ibert_7series_gtp_3750
(
  // GT top level ports
  output [(4*`C_NUM_QUADS)-1:0]		TXN_O,
  output [(4*`C_NUM_QUADS)-1:0]		TXP_O,
  input  [(4*`C_NUM_QUADS)-1:0]    	RXN_I,
  input  [(4*`C_NUM_QUADS)-1:0]   	RXP_I,
  input                           	SYSCLKP_I,
  input  [`C_REFCLKS_USED-1:0]     	GTREFCLK0P_I,
  input  [`C_REFCLKS_USED-1:0]     	GTREFCLK0N_I,
  input  [`C_REFCLKS_USED-1:0]     	GTREFCLK1P_I,
  input  [`C_REFCLKS_USED-1:0]    	GTREFCLK1N_I,
  output                           	LA01_P,
  output                           	LA01_N
);

  //
  // Ibert refclk internal signals
  //
  wire   [`C_NUM_QUADS-1:0]        	gtrefclk0_i;
  wire   [`C_NUM_QUADS-1:0]        	gtrefclk1_i;
  wire   [`C_REFCLKS_USED-1:0]    	refclk0_i;
  wire   [`C_REFCLKS_USED-1:0]     	refclk1_i;
  wire                            	sysclk_i;
  wire                            	CLKFBOUT;
  wire                            	CLKOUT0;
  

  //
  // Refclk IBUFDS instantiations
  //

    IBUFDS_GTE2 u_buf_q1_clk0
      (
        .O            (refclk0_i[0]),
        .ODIV2        (),
        .CEB          (1'b0),
        .I            (GTREFCLK0P_I[0]),
        .IB           (GTREFCLK0N_I[0])
      );

    IBUFDS_GTE2 u_buf_q1_clk1
      (
        .O            (refclk1_i[0]),
        .ODIV2        (),
        .CEB          (1'b0),
        .I            (GTREFCLK1P_I[0]),
        .IB           (GTREFCLK1N_I[0])
      );

  //
  // Refclk connection from each IBUFDS to respective quads depending on the source selected in gui
  //
  assign gtrefclk0_i[0] = refclk0_i[0];
  assign gtrefclk1_i[0] = refclk1_i[0];



  //
  // Sysclock connection
  //
  assign sysclk_i = SYSCLKP_I;


  PLLE2_BASE #(
     .BANDWIDTH("LOW"),
     .CLKIN1_PERIOD(10.0),
     .CLKFBOUT_MULT(10),
     .CLKOUT0_DIVIDE(8),
     .DIVCLK_DIVIDE(1),
     .REF_JITTER1(0.0)
  )
  PLLE2_BASE_inst (
     .CLKOUT0(CLKOUT0),
     .CLKFBOUT(CLKFBOUT),
     .CLKFBIN(CLKFBOUT),
     .CLKIN1(sysclk_i),
     .PWRDWN(1'b0),
     .RST(1'b0)
  );

   ODDR ODDR_inst_P(
      .Q(LA01_P),
      .C(CLKOUT0),
      .CE(1'b1),
      .D1(1'b1),
      .D2(1'b0),
      .R(1'b0),
      .S(1'b0)
   );

   ODDR ODDR_inst_N (
      .Q(LA01_N),
      .C(CLKOUT0),
      .CE(1'b1),
      .D1(1'b0),
      .D2(1'b1),
      .R(1'b0),
      .S(1'b0)
   );

  //
  // IBERT core instantiation
  //
  ibert_7series_gtp_3750 u_ibert_core
    (
      .TXN_O(TXN_O),
      .TXP_O(TXP_O),
      .RXN_I(RXN_I),
      .RXP_I(RXP_I),
      .SYSCLK_I(sysclk_i),
      .GTREFCLK0_I(gtrefclk0_i),
      .GTREFCLK1_I(gtrefclk1_i)
    );

endmodule
